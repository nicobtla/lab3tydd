library verilog;
use verilog.vl_types.all;
entity adc_vlg_vec_tst is
end adc_vlg_vec_tst;
